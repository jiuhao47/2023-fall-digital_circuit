module ic74hc147(
    input [9:0] i,
    output [3:0] y
);

    reg [3:0] m;
    always @(i)
        casez(i)
        10'b0?????????: m=~(4'd9);
        10'b10????????: m=~(4'd8);
        10'b110???????: m=~(4'd7);
        10'b1110??????: m=~(4'd6);
        10'b11110?????: m=~(4'd5);
        10'b111110????: m=~(4'd4);
        10'b1111110???: m=~(4'd3);
        10'b11111110??: m=~(4'd2);
        10'b111111110?: m=~(4'd1);
        default: m=~(4'd0);   
        endcase
    assign y=m;
endmodule

//优先编码器
//输出y低有效